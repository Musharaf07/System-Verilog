// SV Event
//Event is triggered before waiting for Event trigger using wait()
module event_exmpl;
  event ev1;
  
  task process1();
    $display("%0t, Before Capturing event",$time);
    #10;
    wait(ev1.triggered);
    $display("%0t, After Capturing event",$time);
  endtask
  
  task process2();
    $display("%0t, Before triggering event",$time);
    
    #5;
    ->ev1;
    $display("%0t, After triggering event",$time);
 endtask

  initial begin
    fork
      process1();
      process2();
    join
  end
  
endmodule
